module fv_fifo#(

);



/////// Assumptionss//////////////////////
  

/////// Assertions //////////////////////
   
   
/////// Cover properties/////////////////
        


endmodule


bind fifo fv_fifo fv_fifo_inst(.*);
