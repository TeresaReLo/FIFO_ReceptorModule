module fifo_receptor #(
  	
);

  	
 
endmodule

